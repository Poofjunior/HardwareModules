module TickTimeToVelocityLookup(
/// TODO: figure out bit width of input time_per_tick.
            input logic [13:0] time_per_tick,
/// TODO: figure out bit width of output velocity value.
           output logic [15:0] velocity);


endmodule
