`define HARDWARE_MODULES_DIR(filepath) `"/home/poofjunior/Projects/HardwareModules/filepath`" 

